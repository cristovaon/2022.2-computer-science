// Write your modules here!
parameter NUM_OF_BITS=8
module fullAdder(
  input logic signed [NUM_OF_BITS-1:0] number1, number2
  output logic [NUM_OF_BITS-1:0] S);
  
  always_comb begin
  S = A+B
  end
  
  
endmodule
