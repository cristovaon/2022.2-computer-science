/*
Problema 01 - Irrigação
Cristovão Pessoa Cândido Neto - 121110199
*/
module circuit(
  input logic[1:0] U,
  output logic[1:0] S
);
always_comb S <= U;
endmodule
